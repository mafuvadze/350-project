module vga_controller3();


endmodule