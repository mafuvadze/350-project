//// megafunction wizard: %ROM: 1-PORT%VBB%
//// GENERATION: STANDARD
//// VERSION: WM1.0
//// MODULE: altsyncram 
//
//// ============================================================
//// File Name: imem.v
//// Megafunction Name(s):
//// 			altsyncram
////
//// Simulation Library Files(s):
//// 			altera_mf
//// ============================================================
//// ************************************************************
//// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
////
//// 17.1.0 Build 590 10/25/2017 SJ Lite Edition
//// ************************************************************
//
////Copyright (C) 2017  Intel Corporation. All rights reserved.
////Your use of Intel Corporation's design tools, logic functions 
////and other software and tools, and its AMPP partner logic 
////functions, and any output files from any of the foregoing 
////(including device programming or simulation files), and any 
////associated documentation or information are expressly subject 
////to the terms and conditions of the Intel Program License 
////Subscription Agreement, the Intel Quartus Prime License Agreement,
////the Intel FPGA IP License Agreement, or other applicable license
////agreement, including, without limitation, that your use is for
////the sole purpose of programming logic devices manufactured by
////Intel and sold by Intel or its authorized distributors.  Please
////refer to the applicable agreement for further details.
//
//module imem (
//	address,
//	clock,
//	q);
//
//	input	[11:0]  address;
//	input	  clock;
//	output	[31:0]  q;
//`ifndef ALTERA_RESERVED_QIS
//// synopsys translate_off
//`endif
//	tri1	  clock;
//`ifndef ALTERA_RESERVED_QIS
//// synopsys translate_on
//`endif
//
//endmodule
//
//// ============================================================
//// CNX file retrieval info
//// ============================================================
//// Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
//// Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
//// Retrieval info: PRIVATE: AclrByte NUMERIC "0"
//// Retrieval info: PRIVATE: AclrOutput NUMERIC "0"
//// Retrieval info: PRIVATE: BYTE_ENABLE NUMERIC "0"
//// Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
//// Retrieval info: PRIVATE: BlankMemory NUMERIC "0"
//// Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
//// Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
//// Retrieval info: PRIVATE: Clken NUMERIC "0"
//// Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
//// Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
//// Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
//// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
//// Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
//// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
//// Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
//// Retrieval info: PRIVATE: MIFfilename STRING "imem.mif"
//// Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "4096"
//// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
//// Retrieval info: PRIVATE: RegAddr NUMERIC "1"
//// Retrieval info: PRIVATE: RegOutput NUMERIC "1"
//// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
//// Retrieval info: PRIVATE: SingleClock NUMERIC "1"
//// Retrieval info: PRIVATE: UseDQRAM NUMERIC "0"
//// Retrieval info: PRIVATE: WidthAddr NUMERIC "12"
//// Retrieval info: PRIVATE: WidthData NUMERIC "32"
//// Retrieval info: PRIVATE: rden NUMERIC "0"
//// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
//// Retrieval info: CONSTANT: ADDRESS_ACLR_A STRING "NONE"
//// Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
//// Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
//// Retrieval info: CONSTANT: INIT_FILE STRING "imem.mif"
//// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
//// Retrieval info: CONSTANT: LPM_HINT STRING "ENABLE_RUNTIME_MOD=NO"
//// Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
//// Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "4096"
//// Retrieval info: CONSTANT: OPERATION_MODE STRING "ROM"
//// Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
//// Retrieval info: CONSTANT: OUTDATA_REG_A STRING "CLOCK0"
//// Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "12"
//// Retrieval info: CONSTANT: WIDTH_A NUMERIC "32"
//// Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
//// Retrieval info: USED_PORT: address 0 0 12 0 INPUT NODEFVAL "address[11..0]"
//// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
//// Retrieval info: USED_PORT: q 0 0 32 0 OUTPUT NODEFVAL "q[31..0]"
//// Retrieval info: CONNECT: @address_a 0 0 12 0 address 0 0 12 0
//// Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
//// Retrieval info: CONNECT: q 0 0 32 0 @q_a 0 0 32 0
//// Retrieval info: GEN_FILE: TYPE_NORMAL imem.v TRUE
//// Retrieval info: GEN_FILE: TYPE_NORMAL imem.inc FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL imem.cmp FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL imem.bsf FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL imem_inst.v FALSE
//// Retrieval info: GEN_FILE: TYPE_NORMAL imem_bb.v TRUE
//// Retrieval info: LIB_FILE: altera_mf
